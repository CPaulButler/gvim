-------------------------------------------------------------------------------
--
-- File: PkgNewPackage.vhd
-- Author: Paul Butler
-- Original Project: PkgNewPackage
-- Date: TodaysDate
--
-------------------------------------------------------------------------------
-- (c) ThisYear Copyright National Instruments Corporation
-- All Rights Reserved
-- National Instruments Internal Information
-------------------------------------------------------------------------------
--
-- Purpose:
--

library IEEE;
  use IEEE.std_logic_1164.all;

library WORK;
  use WORK.PkgNiUtilities.all;

package PkgNewPackage is
end package PkgNewPackage;

-- The package body is unnecessary if the package contains no subprogram 
-- declarations.
--package body PkgNewPackage is
--end package body PkgNewPackage;

